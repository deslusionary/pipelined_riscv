///////////////////////////////////////////////
// Filename:  reg_file.sv
// Author: Christopher Tinker
// Date: 2022-01-30
//
// Description:
// 	2 read port, 1 write port register file for an
// in-order RV32 processor. Asynchronous read, 
// synchronous (negedge triggered) write.
///////////////////////////////////////////////


module reg_file (

    );
    
endmodule
